library ieee;
use ieee.std_logic_1164.all;
use work.sim_avalon.all;
use ieee.numeric_std.all;
-------------------------------------------------------------------------------

entity mm_bus_seven_seg_four_digit_tb is

end mm_bus_seven_seg_four_digit_tb;

-------------------------------------------------------------------------------

architecture tb of mm_bus_seven_seg_four_digit_tb is
--package sim_avalon is

--  procedure avalon_mm_write (
--    constant write_wait_time : in  integer;
--    constant wr_addr         : in  std_logic_vector(7 downto 0);
--    constant wr_data         : in  std_logic_vector(15 downto 0);
--    signal avs_s1_clk        : in  std_logic;
--    signal avs_s1_cs         : out std_logic;
--    signal avs_s1_write      : out std_logic;
--    signal avs_s1_address    : out std_logic_vector(7 downto 0);
--    signal avs_s1_writedata  : out std_logic_vector(15 downto 0));
--
--  procedure avalon_mm_read (
--    constant read_wait_time : in  integer;
--    constant rd_addr        : in  std_logic_vector(7 downto 0);
--    signal avs_s1_clk       : in  std_logic;
--    signal avs_s1_cs        : out std_logic;
--    signal avs_s1_read      : out std_logic;
--    signal avs_s1_address   : out std_logic_vector(7 downto 0);
--    signal avs_s1_readdata  : in  std_logic_vector(15 downto 0));
--avalon_mm_read(0,"0000000",avs_s1_clk, avs_s1_cs, avs_s1_read, avs_s1_address, avs_s1_readdata);
--end sim_avalon;
function bin27seg (bin : unsigned(3 downto 0)) return std_logic_vector is
variable hex : std_logic_vector(6 downto 0);
begin
   case bin is
      when "0000" => hex := "1000000";  -- 0
      when "0001" => hex := "1111001";  -- 1
      when "0010" => hex := "0100100";  -- 2
      when "0011" => hex := "0110000";  -- 3
      when "0100" => hex := "0011001";  -- 4
      when "0101" => hex := "0010010";  -- 5
      when "0110" => hex := "0000010";  -- 6
      when "0111" => hex := "1111000";  -- 7
      when "1000" => hex := "0000000";  -- 8
      when "1001" => hex := "0011000";  -- 9
      when "1010" => hex := "0001000";  -- a
      when "1011" => hex := "0000011";  -- b
      when "1100" => hex := "1000110";  -- c
      when "1101" => hex := "0100001";  -- d
      when "1110" => hex := "0000110";  -- e
      when "1111" => hex := "0001110";  -- f
      when others => null;
    end case;
    return hex;
end bin27seg;

  component mm_bus_seven_seg_four_digit
    port (
      csi_clockreset_clk     : in  std_logic;
      csi_clockreset_reset_n : in  std_logic;
      avs_s1_write           : in  std_logic;
      avs_s1_read            : in  std_logic;
      avs_s1_chipselect      : in  std_logic;
      avs_s1_address         : in  std_logic_vector(7 downto 0);
      avs_s1_writedata       : in  std_logic_vector(15 downto 0);
      avs_s1_readdata        : out std_logic_vector(15 downto 0);
      hex0                   : out std_logic_vector(6 downto 0);
      hex1                   : out std_logic_vector(6 downto 0);
      hex2                   : out std_logic_vector(6 downto 0);
      hex3                   : out std_logic_vector(6 downto 0));
  end component;

  -- constants
  constant read_wait_time  : integer := 1;
  constant write_wait_time : integer := 2;

  -- component ports
  signal csi_clockreset_clk     : std_logic := '0';
  signal csi_clockreset_reset_n : std_logic := '1';
  signal avs_s1_write           : std_logic := '0';
  signal avs_s1_read            : std_logic := '0';
  signal avs_s1_chipselect      : std_logic := '0';
  signal avs_s1_address         : std_logic_vector(7 downto 0) := (others => '0');
  signal avs_s1_writedata       : std_logic_vector(15 downto 0) := (others => '0');
  signal avs_s1_readdata        : std_logic_vector(15 downto 0) := (others => 'Z');
  signal hex0                   : std_logic_vector(6 downto 0) := (others => '1');
  signal hex1                   : std_logic_vector(6 downto 0) := (others => '1');
  signal hex2                   : std_logic_vector(6 downto 0) := (others => '1');
  signal hex3                   : std_logic_vector(6 downto 0) := (others => '1');

  -- clock
  signal Clk : std_logic := '1';
	signal running : std_logic := '1';
begin  -- tb

  -- component instantiation
  DUT: mm_bus_seven_seg_four_digit
    port map (
      csi_clockreset_clk     => csi_clockreset_clk,
      csi_clockreset_reset_n => csi_clockreset_reset_n,
      avs_s1_write           => avs_s1_write,
      avs_s1_read            => avs_s1_read,
      avs_s1_chipselect      => avs_s1_chipselect,
      avs_s1_address         => avs_s1_address,
      avs_s1_writedata       => avs_s1_writedata,
      avs_s1_readdata        => avs_s1_readdata,
      hex0                   => hex0,
      hex1                   => hex1,
      hex2                   => hex2,
      hex3                   => hex3);

  -- clock generation
  
  Clk <= not Clk after 10 ns;
  csi_clockreset_clk <= Clk;
  csi_clockreset_reset_n <= '0', '1' after 5 ns;

  -- waveform generation
  WaveGen_Proc: process
  variable bin : unsigned(15 downto 0);
  variable hex_tmp : std_logic_vector(6 downto 0);
  begin
	
	wait until csi_clockreset_clk = '0';
	wait until csi_clockreset_clk = '1';
	bin(15 downto 12) := to_unsigned(1,4);
	bin(11 downto 8) := to_unsigned(2,4);
	bin(7 downto 4) := to_unsigned(3,4);
	bin(3 downto 0) := to_unsigned(4,4);
	avalon_mm_write(1,"00000000",std_logic_vector(bin),csi_clockreset_clk, avs_s1_chipselect, avs_s1_write, avs_s1_address, avs_s1_writedata);
	
	wait until csi_clockreset_clk = '0';
	wait until csi_clockreset_clk = '1';
	--hex_tmp := bin27seg(bin(3 downto 0)) ;
	assert hex0 = bin27seg(bin(3 downto 0))
		and hex1 = bin27seg(bin(7 downto 4))
		and hex2 = bin27seg(bin(11 downto 8)) 
		and hex3 = bin27seg(bin(15 downto 12))
			report "7seg driver not working!!"
				severity failure;
	report "done"
		severity note;
    wait;
  end process WaveGen_Proc;

end tb;

-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
